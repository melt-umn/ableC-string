grammar edu:umn:cs:melt:exts:ableC:string;

exports edu:umn:cs:melt:exts:ableC:string:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:string:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:templating;
